
	/*==========================================================*/

    /*generate ten data and one data

	/*==========================================================*/
	





    /***********************************************************/





    /*==========================================================*/
